package fifo_env_pkg;

import uvm_pkg::*;
import fifo_stimulus_pkg::*;

`include "fifo_driver.sv"
`include "fifo_monitor.sv"
`include "fifo_agent.sv"
`include "fifo_scoreboard.sv"
`include "fifo_env.sv"

endpackage: fifo_env_pkg
