package fifo_test_pkg;

import uvm_pkg::*;
import fifo_stimulus_pkg::*;
import fifo_env_pkg::*;

`include "test_collection.sv"

endpackage: fifo_test_pkg
