package fifo_stimulus_pkg;

import uvm_pkg::*;
`include "fifo_item.sv"
`include "fifo_item_ow.sv"
`include "fifo_sequence.sv"

endpackage: fifo_stimulus_pkg
